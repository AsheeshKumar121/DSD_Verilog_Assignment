`timescale 1ns / 1ps

module OR_Design(
input a,
input b,
output y
    );
    
    assign y=a|b;
    
endmodule