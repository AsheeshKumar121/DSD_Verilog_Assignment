`timescale 1ns / 1ps

module NOT_Design(
input a,
output y
    );
    
    assign y = ~a;
    
endmodule