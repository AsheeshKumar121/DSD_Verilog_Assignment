`timescale 1ns / 1ps

module XNOR_Design(
input a,b,
output y
    );
    
    assign y = ~(a^b);
    
endmodule